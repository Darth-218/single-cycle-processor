module alu_contorl_test;
endmodule
