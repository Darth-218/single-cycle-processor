module single_cycle_processor_test;
endmodule

