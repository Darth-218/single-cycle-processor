module alu_control_test;
endmodule
